
.subckt TOP
C1 A B 1f
.ends

