
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPD0 y D1 pndC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMND0 y D1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPD0 y D1 pndC VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 y D1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPD0 y D1 pndC VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMND0 y D1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPD0 Y D1 pndC VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 Y D1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPD0 Y D1 pndC VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 Y D1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPC0 pndC C1 pndB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPD0 Y D1 pndC VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMND0 Y D1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a2111oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a211oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21bo_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21bo_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21bo_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 net40 A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 net40 A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 net40 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__a21boi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 net40 A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 net40 A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 net40 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__a21boi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 net40 A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 net40 A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 net40 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21boi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a21oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a221oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 y C2 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 net68 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI10 net68 C2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__a222o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a222o_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI8 y C2 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 net68 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI10 net68 C2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__a222o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MI8 Y C2 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 Y C1 net62 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI10 net62 C2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__a222oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a222oi_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 pndB B2 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MI8 Y C2 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 Y C1 net62 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI10 net62 C2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__a222oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a22oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi11 sndNB1 B2 y VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi20 y inor VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMPaoi20 y inor pmid VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 sndNB1 B2 y VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 y inor VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPaoi20 y inor pmid VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi11 sndNB1 B2 y VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi20 y inor VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPaoi20 y inor pmid VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 Y inor VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi20 Y inor pmid VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi20 Y inor VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi20 Y inor pmid VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnor0 inor A1_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnor1 inor A2_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi20 Y inor VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPaoi10 pmid B1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi11 pmid B2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi20 Y inor pmid VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__a2bb2oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 y C1 pndB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 pndB B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPC0 Y C1 pndB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a311oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a31oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 y B2 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 Y B2 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 sndA2 A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 sndB1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 sndB1 B2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a32oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41o_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41o_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 y B1 pndA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41o_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41oi_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41oi_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 pndA A1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 pndA A2 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 pndA A3 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA3 pndA A4 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 Y B1 pndA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 Y A1 sndA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA3 sndA3 A4 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__a41oi_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2b_1 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2b_2 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and2b_4 A_N B VGND VNB VPB VPWR X
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3b_1 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3b_2 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and3b_4 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and3b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4_1 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4_2 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4_4 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4b_1 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4b_2 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4b_4 A_N B C D VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4bb_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4bb_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 y C VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 y D VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and4bb_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__buf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__buf_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=6 w=0.74 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=16 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=6 w=1.12 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=16 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__buf_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__buf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__buf_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__buf_4 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__buf_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__buf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=3 w=0.74 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=8 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__buf_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__bufbuf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 Abb Ab VGND VNB nfet_01v8_lvt m=3 w=0.74 l=0.15
MMIN3 Abbb Abb VGND VNB nfet_01v8_lvt m=6 w=0.74 l=0.15
MMIN4 X Abbb VGND VNB nfet_01v8_lvt m=16 w=0.74 l=0.15
MMIP4 X Abbb VPWR VPB pfet_01v8 m=16 w=1.12 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP2 Abb Ab VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
MI5 Abbb Abb VPWR VPB pfet_01v8 m=6 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__bufbuf_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__bufbuf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 Abbb Abb VGND VNB nfet_01v8_lvt m=3 w=0.74 l=0.15
MMIN4 X Abbb VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIP4 X Abbb VPWR VPB pfet_01v8 m=8 w=1.12 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI5 Abbb Abb VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__bufbuf_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__bufinv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=3 w=0.74 l=0.15
MMIN2 Abb Ab VGND VNB nfet_01v8_lvt m=6 w=0.74 l=0.15
MMIN3 Y Abb VGND VNB nfet_01v8_lvt m=16 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
MMIP2 Abb Ab VPWR VPB pfet_01v8 m=6 w=1.12 l=0.15
MMIP3 Y Abb VPWR VPB pfet_01v8 m=16 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__bufinv_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__bufinv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 Abb Ab VGND VNB nfet_01v8_lvt m=3 w=0.74 l=0.15
MMIN3 Y Abb VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIP1 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP2 Abb Ab VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
MMIP3 Y Abb VPWR VPB pfet_01v8 m=8 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__bufinv_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN0 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN1 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP0 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkbuf_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN0 Ab A VGND VNB nfet_01v8_lvt m=4 w=0.42 l=0.15
MMIN1 X Ab VGND VNB nfet_01v8_lvt m=16 w=0.42 l=0.15
MMIP0 Ab A VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 X Ab VPWR VPB pfet_01v8 m=16 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkbuf_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkbuf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN0 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN1 X Ab VGND VNB nfet_01v8_lvt m=2 w=0.42 l=0.15
MMIP0 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 X Ab VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkbuf_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkbuf_4 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN0 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN1 X Ab VGND VNB nfet_01v8_lvt m=4 w=0.42 l=0.15
MMIP0 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 X Ab VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkbuf_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkbuf_8 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN0 Ab A VGND VNB nfet_01v8_lvt m=2 w=0.42 l=0.15
MMIN1 X Ab VGND VNB nfet_01v8_lvt m=8 w=0.42 l=0.15
MMIP0 Ab A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 X Ab VPWR VPB pfet_01v8 m=8 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkbuf_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv3sd1_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 Y Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1 l=0.15
MMIP2 Y Abb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkdlyinv3sd1_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv3sd2_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 Y Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1 l=0.25
MMIP2 Y Abb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkdlyinv3sd2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv3sd3_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 Y Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.5
MMIP2 Y Abb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkdlyinv3sd3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv5sd1_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 Y Abbbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 Abbbb Abbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI13 Abbb Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 Y Abbbb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 Abbbb Abbb VPWR VPB pfet_01v8 m=1 w=1 l=0.15
MI14 Abbb Abb VPWR VPB pfet_01v8 m=1 w=1 l=0.15
.ENDS sky130_fd_sc_hs__clkdlyinv5sd1_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv5sd2_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 Y Abbbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 Abbbb Abbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MI13 Abbb Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.25
MMIP2 Y Abbbb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 Abbbb Abbb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.25
MI14 Abbb Abb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.25
.ENDS sky130_fd_sc_hs__clkdlyinv5sd2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkdlyinv5sd3_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 Y Abbbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 Abbbb Abbb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MI13 Abbb Abb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIP1 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.5
MMIP2 Y Abbbb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 Abbbb Abbb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.5
MI14 Abbb Abb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.5
.ENDS sky130_fd_sc_hs__clkdlyinv5sd3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkinv_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIP0 Y A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__clkinv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkinv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN0 Y A VGND VNB nfet_01v8_lvt m=16 w=0.42 l=0.15
MMIP0 Y A VPWR VPB pfet_01v8 m=24 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkinv_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkinv_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.42 l=0.15
MMIP0 Y A VPWR VPB pfet_01v8 m=3 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkinv_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkinv_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN0 Y A VGND VNB nfet_01v8_lvt m=4 w=0.42 l=0.15
MMIP0 Y A VPWR VPB pfet_01v8 m=6 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkinv_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__clkinv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN0 Y A VGND VNB nfet_01v8_lvt m=8 w=0.42 l=0.15
MMIP0 Y A VPWR VPB pfet_01v8 m=12 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__clkinv_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__conb_1 VGND VNB VPB VPWR HI LO
*.PININFO VGND:I VNB:I VPB:I VPWR:I HI:O LO:O
*rI12 VGND LO short
*rI11 HI VPWR short
.ENDS sky130_fd_sc_hs__conb_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__decap_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
MI2 VPWR VGND VPWR VPB pfet_01v8 m=1 w=1.0 l=1.0
MI1 VGND VPWR VGND VNB nfet_01v8_lvt m=1 w=0.42 l=1.0
.ENDS sky130_fd_sc_hs__decap_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI659 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net141 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net162 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI677 M1 RESET net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net125 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net125 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 net82 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net82 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 net162 net82 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net93 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net93 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net82 RESET net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net82 S0 net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net81 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net218 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net162 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI9 net82 S0 net221 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net218 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net165 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net210 net82 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net210 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net82 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net221 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net194 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI665 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI656 M0 clkneg net194 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net165 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net162 net82 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI661 Q_N net82 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfbbn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI659 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net141 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net162 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI677 M1 RESET net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net118 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net118 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 net82 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net82 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI652 net162 net82 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net93 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net93 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net82 RESET net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net82 S0 net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net81 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net218 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net162 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI9 net82 S0 net221 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net218 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net165 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net210 net82 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net210 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net82 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net221 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net194 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI665 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI656 M0 clkneg net194 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net165 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net162 net82 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI661 Q_N net82 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfbbn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI659 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net141 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net162 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI677 M1 RESET net141 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net125 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net125 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 net82 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net82 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 net162 net82 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net93 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net93 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net82 RESET net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net82 S0 net81 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net81 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net218 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net162 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI9 net82 S0 net221 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net218 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net165 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net210 net82 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net210 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net82 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net221 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net194 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI665 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI656 M0 clkneg net194 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net165 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net162 net82 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI661 Q_N net82 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfbbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI651 Q_N s0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net93 s0 net123 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net123 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net116 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net108 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net108 M1 net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net92 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net168 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net168 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net92 net93 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI39 db D net76 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net76 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net196 net93 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net93 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net196 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net93 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net175 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net175 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net168 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net168 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI661 Q_N s0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI651 Q_N s0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net93 s0 net123 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net123 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net116 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net108 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net108 M1 net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net92 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net168 s0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI653 Q net168 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI654 net92 net93 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D net76 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net76 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net196 net93 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net93 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net196 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net93 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net175 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net175 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net168 s0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net168 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI661 Q_N s0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK_N:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net88 s0 net118 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net118 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net111 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net103 M1 net111 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net87 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net155 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net155 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net87 net88 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net71 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net183 net88 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net88 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net183 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net88 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net162 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net162 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net155 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net155 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrtn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net88 s0 net118 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net118 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net111 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net103 M1 net111 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net87 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net155 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net155 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net87 net88 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net71 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net183 net88 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net88 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net183 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net88 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net162 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net162 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net155 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net155 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net88 s0 net118 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net118 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net111 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net103 M1 net111 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net87 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net155 s0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 Q net155 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI654 net87 net88 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net71 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net183 net88 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net88 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net183 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net88 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net162 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net162 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net155 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net155 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net88 s0 net118 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net118 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net111 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net103 M1 net111 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net87 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net155 s0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 Q net155 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI654 net87 net88 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI38 net71 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net183 net88 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net88 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net183 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net88 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net162 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net162 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net155 s0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI660 Q net155 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI41 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__dfrtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI36 net129 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net112 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net80 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net129 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI25 net97 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI26 S0 clkneg net89 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net89 S1 net97 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net80 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net112 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net141 S0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net141 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI49 Q_N S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net192 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net192 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net169 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net169 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net156 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI5 S0 clkpos net156 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net141 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net141 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI50 Q_N S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfsbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI36 net128 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net111 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net108 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net128 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI25 net96 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI26 S0 clkneg net88 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net88 S1 net96 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net108 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net111 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net140 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI653 Q net140 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI49 Q_N S0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net191 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net191 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net168 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net168 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net155 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI5 S0 clkpos net155 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net140 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net140 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI50 Q_N S0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfsbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI36 net120 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net71 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net120 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI25 net88 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI26 S0 clkneg net80 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net80 S1 net88 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net103 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net128 S0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net128 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net179 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net179 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net156 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net156 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net143 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI5 S0 clkpos net143 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net128 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net128 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfstp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI36 net120 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net71 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net120 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI25 net88 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI26 S0 clkneg net80 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net80 S1 net88 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net103 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net128 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI653 Q net128 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net179 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net179 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net156 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net156 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net143 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI5 S0 clkpos net143 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net128 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net128 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfstp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI36 net120 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI39 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net103 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net71 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net120 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI25 net88 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI26 S0 clkneg net80 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net80 S1 net88 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net103 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net128 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 Q net128 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI40 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net179 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net179 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net156 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net156 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net143 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI5 S0 clkpos net143 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net128 S0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI660 Q net128 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfstp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI657 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net96 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI669 net88 S1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net72 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net72 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI665 Q_N net88 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI659 M0 clkneg net128 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI644 S0 clkpos net147 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI670 net88 S1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI643 net147 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net128 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI666 Q_N net88 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfxbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI657 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net96 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net76 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net76 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI669 net52 S1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI665 Q_N net52 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI659 M0 clkneg net132 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI644 S0 clkpos net147 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI643 net147 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net132 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI670 net52 S1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI666 Q_N net52 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfxbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI657 M0 clkpos net79 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net79 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net59 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net59 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI659 M0 clkneg net107 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net122 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI643 net122 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net107 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfxtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfxtp_2 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI657 M0 clkpos net79 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net79 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net59 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net59 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI659 M0 clkneg net107 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI644 S0 clkpos net122 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI643 net122 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net107 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfxtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI657 M0 clkpos net79 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net79 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 db D VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net59 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net59 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI659 M0 clkneg net107 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI644 S0 clkpos net122 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI643 net122 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net107 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 db D VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__dfxtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__diode_2 DIODE VGND VNB VPB VPWR
*.PININFO DIODE:I VGND:I VNB:I VPB:I VPWR:I
* Notes: Tap diode is not represented here.
.ENDS sky130_fd_sc_hs__diode_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net75 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net75 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net63 CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 net63 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI38 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net54 GATE VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net63 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 M0 clkpos net91 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net99 CLK VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI656 net63 m1 net99 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI36 net91 GATE VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net63 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__dlclkp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net75 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net75 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net63 CLK VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI658 net63 m1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI38 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net54 GATE VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net63 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 M0 clkpos net91 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net99 CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net63 m1 net99 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI36 net91 GATE VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net63 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__dlclkp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net75 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net75 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net63 CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net63 m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI38 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net54 GATE VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net63 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net110 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net110 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 M0 clkpos net91 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net99 CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net63 m1 net99 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI36 net91 GATE VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net63 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__dlclkp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net125 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 M0 clkneg net61 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net125 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net61 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net57 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net57 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net125 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI645 net125 m1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net116 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net121 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net96 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrbn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net125 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI17 M0 clkneg net61 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net125 m1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net61 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net57 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net57 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net125 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI645 net125 m1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net108 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net116 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net108 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net96 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrbn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net125 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 M0 clkneg net61 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net125 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net61 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net57 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net57 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net125 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI645 net125 m1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net116 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net121 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net96 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net125 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI17 M0 clkneg net61 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net125 m1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net61 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net57 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net57 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net125 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI645 net125 m1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net108 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net116 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net116 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net108 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net96 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net96 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI18 net54 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net50 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net50 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net106 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net101 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net101 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net106 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net81 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net81 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net54 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net50 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net50 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI657 net106 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net101 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net101 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net106 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net81 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net81 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net55 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI18 net55 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net51 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net51 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI657 net94 RESET_B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI652 M0 clkneg net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net102 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net94 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net82 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net82 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtn_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI18 net54 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net50 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net50 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net93 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net101 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net101 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net93 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net81 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net81 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net54 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI18 net54 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net50 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net50 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI657 net93 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net101 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net101 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net93 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net81 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net81 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I RESET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net55 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 m1 RESET_B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI18 net55 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net51 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net51 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI657 net94 RESET_B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI652 M0 clkneg net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net102 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 net94 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net82 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net82 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlrtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net112 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 M0 clkneg net56 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net112 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net56 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net52 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net52 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net112 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI645 net112 m1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI652 M0 clkneg net107 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net107 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net87 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net87 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxbn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net114 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI17 M0 clkneg net58 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net114 m1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net58 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net54 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net54 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net114 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI645 net114 m1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI652 M0 clkneg net109 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net109 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net89 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net89 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxbn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
*.PININFO D:I GATE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI648 Q_N net114 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 M0 clkneg net58 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI646 net114 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net58 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net54 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net54 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI647 Q_N net114 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI645 net114 m1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI652 M0 clkneg net109 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net109 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net89 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net89 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net53 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net53 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net44 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net44 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net96 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net96 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net76 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net76 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxtn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net51 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net51 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net47 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net47 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI652 M0 clkneg net94 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net94 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net74 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net74 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxtn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
*.PININFO D:I GATE_N:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net51 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI633 clkpos GATE_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net51 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net47 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net47 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkpos GATE_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI652 M0 clkneg net94 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net94 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net74 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 net74 db VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__dlxtn_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlxtp_1 D GATE VGND VNB VPB VPWR Q
*.PININFO D:I GATE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI17 M0 clkneg net51 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 Q m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI633 clkneg GATE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI18 net51 db VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI653 net47 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 M0 clkpos net47 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI655 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI638 db D VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI634 clkneg GATE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 Q m1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 M0 clkneg net94 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net94 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI637 db D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI19 M0 clkpos net74 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI20 net74 db VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__dlxtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlygate4sd1_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab net34 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net34 net30 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 net30 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Ab net34 VPWR VPB pfet_01v8 m=1 w=1 l=0.18
MMIP2 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 net34 net30 VPWR VPB pfet_01v8 m=1 w=1 l=0.18
MI8 net30 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlygate4sd1_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlygate4sd2_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab net34 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net34 net30 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MI9 net30 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Ab net34 VPWR VPB pfet_01v8 m=1 w=1 l=0.25
MMIP2 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 net34 net30 VPWR VPB pfet_01v8 m=1 w=1 l=0.25
MI8 net30 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlygate4sd2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlygate4sd3_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab net34 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net34 net30 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.18
MI9 net30 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIP1 Ab net34 VPWR VPB pfet_01v8 m=1 w=1 l=0.5
MMIP2 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 net34 net30 VPWR VPB pfet_01v8 m=1 w=1 l=0.5
MI8 net30 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlygate4sd3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlymetal6s2s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab net055 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 net47 Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net055 net59 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI15 net55 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 net59 X VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 X net55 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP1 Ab net055 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MMIP2 net47 Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 net055 net59 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 net59 X VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI18 X net55 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 net55 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlymetal6s2s_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlymetal6s4s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab X VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 net47 Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 X net59 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI15 net55 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 net59 net63 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net63 net55 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP1 Ab X VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MMIP2 net47 Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 X net59 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 net59 net63 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI18 net63 net55 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 net55 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlymetal6s4s_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__dlymetal6s6s_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab net055 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMIN2 X Ab VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net055 net59 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI15 net55 A VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI9 net59 net63 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net63 net55 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP1 Ab net055 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MMIP2 X Ab VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI7 net055 net59 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI8 net59 net63 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI18 net63 net55 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI17 net55 A VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__dlymetal6s6s_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ebufn_1 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z net35 sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA net39 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 net39 TE_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI6 net35 A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndTEB net35 Z VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 net39 TE_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI5 net35 A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__ebufn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ebufn_2 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z net35 sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA net39 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 net39 TE_B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI6 net35 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndTEB net35 Z VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 net39 TE_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI5 net35 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__ebufn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ebufn_4 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z net35 sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA net39 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN1 net39 TE_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net35 A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndTEB net35 Z VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 net39 TE_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI5 net35 A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__ebufn_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ebufn_8 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z net35 sndA VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMN1 sndA net39 VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIN1 net39 TE_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 net35 A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=8 w=1.12 l=0.15
MMP1 sndTEB net35 Z VPB pfet_01v8 m=8 w=1.12 l=0.15
MMIP1 net39 TE_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI5 net35 A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__ebufn_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI14 net123 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net123 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI655 net63 deneg VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net108 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net91 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net91 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI660 Q_N S1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M0 clkneg net108 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net80 DE VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI9 db S1 net80 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI4 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI8 db D net63 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI661 Q_N S1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net188 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net188 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net143 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net163 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net163 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI16 net156 M1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI15 S0 clkpos net156 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI5 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI7 db D net143 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI11 db S1 net136 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI12 net136 deneg VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__edfxbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI14 net115 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net115 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI655 net59 deneg VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net79 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net83 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net83 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 M0 clkneg net79 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net76 DE VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI9 db S1 net76 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI4 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI8 db D net59 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net175 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net175 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net172 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net160 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net160 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net148 M1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI15 S0 clkpos net148 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI5 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI7 db D net172 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI11 db S1 net128 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI12 net128 deneg VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__edfxtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvn_1 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA net25 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 net25 TE_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 net25 TE_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__einvn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvn_2 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 TE TE_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 TE TE_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__einvn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvn_4 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN1 TE TE_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 TE TE_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__einvn_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvn_8 A TE_B VGND VNB VPB VPWR Z
*.PININFO A:I TE_B:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIN1 TE TE_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMP0 VPWR TE_B sndTEB VPB pfet_01v8 m=8 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=8 w=1.12 l=0.15
MMIP1 TE TE_B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__einvn_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvp_1 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 TEB TE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMP0 VPWR TEB sndTEB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 TEB TE VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__einvp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvp_2 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 TEB TE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MMP0 VPWR TEB sndTEB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 TEB TE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__einvp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvp_4 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN1 TEB TE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMP0 VPWR TEB sndTEB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 TEB TE VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__einvp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__einvp_8 A TE VGND VNB VPB VPWR Z
*.PININFO A:I TE:I VGND:I VNB:I VPB:I VPWR:I Z:O
MMN0 Z A sndA VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMN1 sndA TE VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIN1 TEB TE VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMP0 VPWR TEB sndTEB VPB pfet_01v8 m=8 w=1.12 l=0.15
MMP1 sndTEB A Z VPB pfet_01v8 m=8 w=1.12 l=0.15
MMIP1 TEB TE VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__einvp_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMNs1s nint1 majb sumb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj10 majb B sndNAp1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs3s0 nint1 B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs3s1 nint1 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs3s2 nint1 CIN VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj11 sndPAp1 B majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s0 pint1 B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s1 pint1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1s pint1 majb sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__fa_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMNs1s nint1 majb sumb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNmaj10 majb B sndNAp1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj30 majb CIN nmajmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj21 nmajmid A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj20 VGND B nmajmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s0 nint1 A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s1 nint1 B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s2 nint1 CIN VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj11 sndPAp1 B majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj20 VPWR B pmajmid VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj30 pmajmid CIN majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj21 pmajmid A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s0 pint1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s1 pint1 B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1s pint1 majb sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__fa_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMNs1s nint1 majb sumb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNmaj10 majb B sndNAp1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj30 majb CIN nmajmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj21 nmajmid A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNmaj20 VGND B nmajmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s0 nint1 A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s1 nint1 B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs3s2 nint1 CIN VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj11 sndPAp1 B majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj20 VPWR B pmajmid VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj30 pmajmid CIN majb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPmaj21 pmajmid A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s0 pint1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s1 pint1 B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1s pint1 majb sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__fa_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT net195 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 SUM net123 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 CIb mid2 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI5 Bb mid1 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 CIbb mid2 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 CIb mid1 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 CIbb CIb VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 CIb CI VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI8 Ab2 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI9 Abb2 Ab2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI14 Ab1 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 Abb2 B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI21 Ab1 Bb mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Abb2 Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Ab1 B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 COUT net195 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP3 SUM net123 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI4 CIb mid1 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI3 Bb mid2 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 CIbb mid1 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 CIb mid2 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 CIbb CIb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI45 CIb CI VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI12 Ab2 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI13 Abb2 Ab2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 Ab1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI22 Abb2 Bb mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI23 Ab1 B mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI26 Abb2 B mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 Ab1 Bb mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__fah_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT net195 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN3 SUM net123 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI6 CIb mid2 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI5 Bb mid1 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 CIbb mid2 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 CIb mid1 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 CIbb CIb VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 CIb CI VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI8 Ab2 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI9 Abb2 Ab2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI14 Ab1 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 Abb2 B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI21 Ab1 Bb mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Abb2 Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Ab1 B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 COUT net195 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP3 SUM net123 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI4 CIb mid1 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI3 Bb mid2 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 CIbb mid1 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 CIb mid2 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 CIbb CIb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI45 CIb CI VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI12 Ab2 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI13 Abb2 Ab2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 Ab1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI22 Abb2 Bb mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI23 Ab1 B mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI26 Abb2 B mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 Ab1 Bb mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__fah_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT net195 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN3 SUM net123 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI6 CIb mid2 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI5 Bb mid1 net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 CIbb mid2 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 CIb mid1 net123 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 CIbb CIb VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 CIb CI VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI8 Ab2 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI9 Abb2 Ab2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI14 Ab1 A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 Abb2 B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI21 Ab1 Bb mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Abb2 Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Ab1 B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 COUT net195 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP3 SUM net123 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI4 CIb mid1 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI3 Bb mid2 net195 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 CIbb mid1 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI650 CIb mid2 net123 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI47 CIbb CIb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI45 CIb CI VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI12 Ab2 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI13 Abb2 Ab2 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 Ab1 A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI22 Abb2 Bb mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI23 Ab1 B mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI26 Abb2 B mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 Ab1 Bb mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__fah_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I CIN:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIP3 SUM net144 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI32 Bbb Bb VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI27 Ab Bb mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI26 Abb B mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI22 Abb Bb mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI23 Ab B mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI19 CINb1 CIN VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI12 CINb2 CIN VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 CINbb2 mid2 net144 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI1 CINb2 mid1 net144 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI3 Bbb mid2 COUT VPB pfet_01v8 m=1 w=0.84 l=0.15
MI4 CINb1 mid1 COUT VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIN3 SUM net144 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 CINb1 mid2 COUT VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Ab B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Abb Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI21 Ab Bb mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 Abb B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI14 CINb1 CIN VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI9 CINbb2 CINb2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI8 CINb2 CIN VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 CINbb2 mid1 net144 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 CINb2 mid2 net144 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI31 Bbb mid1 COUT VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI33 Bbb Bb VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__fahcin_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
*.PININFO A:I B:I CI:I VGND:I VNB:I VPB:I VPWR:I COUT_N:O SUM:O
MMIP3 SUM net146 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI32 Bb2 B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI27 Ab Bb1 mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI26 Abb B mid2 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI22 Abb Bb1 mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI23 Ab B mid1 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI19 CIb1 CI VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI12 CIb2 CI VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI16 Bb1 B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 CIb2 mid2 net146 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI1 CIbb2 mid1 net146 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI3 Bb2 mid2 COUT_N VPB pfet_01v8 m=1 w=0.84 l=0.15
MI4 CIb1 mid1 COUT_N VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIN3 SUM net146 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI6 CIb1 mid2 COUT_N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Ab B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Abb Bb1 mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI21 Ab Bb1 mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI20 Abb B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI14 CIb1 CI VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI9 CIbb2 CIb2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI8 CIb2 CI VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb1 B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 CIb2 mid1 net146 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 CIbb2 mid2 net146 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI31 Bb2 mid1 COUT_N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI33 Bb2 B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__fahcon_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fill_diode_2 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Diffusion diodes are not marked as devices and so not
*        represented here.
.ENDS sky130_fd_sc_hs__fill_diode_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fill_diode_4 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Diffusion diodes are not marked as devices and so not
*        represented here.
.ENDS sky130_fd_sc_hs__fill_diode_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__fill_diode_8 VGND VNB VPB VPWR
*.PININFO VGND:I VNB:I VPB:I VPWR:I
* Notes: Diffusion diodes are not marked as devices and so not
*        represented here.
.ENDS sky130_fd_sc_hs__fill_diode_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ha_1 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA B majb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs1 sumb majb nint1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs20 VGND A nint1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs21 VGND B nint1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPnand0 majb A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 majb B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPs1 VPWR majb sumb VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPs20 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs21 sndPA B sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__ha_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ha_2 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnand1 sndNA B majb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs1 sumb majb nint1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs20 VGND A nint1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs21 VGND B nint1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPnand0 majb A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnand1 majb B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1 VPWR majb sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs20 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs21 sndPA B sumb VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__ha_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__ha_4 A B VGND VNB VPB VPWR COUT SUM
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I COUT:O SUM:O
MMIN2 COUT majb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN3 SUM sumb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNnand1 sndNA B majb VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNs1 sumb majb nint1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNs20 VGND A nint1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNs21 VGND B nint1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIP2 COUT majb VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP3 SUM sumb VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPnand0 majb A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPnand1 majb B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPs1 VPWR majb sumb VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPs20 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPs21 sndPA B sumb VPB pfet_01v8 m=2 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__ha_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__inv_1 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP1 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__inv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Y A VGND VNB nfet_01v8_lvt m=16 w=0.74 l=0.15
MMIP1 Y A VPWR VPB pfet_01v8 m=16 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__inv_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIP1 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__inv_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Y A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIP1 Y A VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__inv_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__inv_8 A VGND VNB VPB VPWR Y
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMIN1 Y A VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMIP1 Y A VPWR VPB pfet_01v8 m=8 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__inv_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__maj3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN10 y B sndNBa VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN11 sndNBa A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN20 y B sndNBc VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN21 sndNBc C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN30 y C sndNCa VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN31 sndNCa A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP10 VPWR A sndPAb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP11 sndPAb B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP20 VPWR C sndPCb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP21 sndPCb B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP30 VPWR A sndPAc VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP31 sndPAc C y VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__maj3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__maj3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN10 y B sndNBa VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN11 sndNBa A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN20 y B sndNBc VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN21 sndNBc C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN30 y C sndNCa VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN31 sndNCa A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP10 VPWR A sndPAb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP11 sndPAb B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP20 VPWR C sndPCb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP21 sndPCb B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP30 VPWR A sndPAc VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP31 sndPAc C y VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__maj3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__maj3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN10 y B sndNBa VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN11 sndNBa A VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN20 y B sndNBc VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN21 sndNBc C VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN30 y C sndNCa VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN31 sndNCa A VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP10 VPWR A sndPAb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP11 sndPAb B y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP20 VPWR C sndPCb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP21 sndPCb B y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP30 VPWR A sndPAc VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP31 sndPAc C y VPB pfet_01v8 m=2 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__maj3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 xb A0 smdNA0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA10 xb A1 sndNA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X xb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA01 sndPS A0 xb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA11 sndPSb A1 xb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X xb VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2_2 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 xb A0 smdNA0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA10 xb A1 sndNA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X xb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA01 sndPS A0 xb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA11 sndPSb A1 xb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X xb VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 xb A0 smdNA0 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA10 xb A1 sndNA1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 X xb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA01 sndPS A0 xb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA11 sndPSb A1 xb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X xb VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNA00 Y A0 smdNA0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA10 Y A1 sndNA1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA01 sndPS A0 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA11 sndPSb A1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__mux2i_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNA00 Y A0 smdNA0 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA10 Y A1 sndNA1 VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA01 sndPS A0 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA11 sndPSb A1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__mux2i_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNA00 Y A0 smdNA0 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA01 smdNA0 Sb VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA10 Y A1 sndNA1 VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA11 sndNA1 S VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN1 Sb S VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPA00 VPWR S sndPS VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA01 sndPS A0 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA10 VPWR Sb sndPSb VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA11 sndPSb A1 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 Sb S VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__mux2i_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs1o xb S1b xlowb VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNs2o xb S1 xhib VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 VGND S1 S1b VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 VGND S0 S0b VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN4 VGND xb X VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1o xb S1 xlowb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2o xb S1b xhib VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 VPWR S1 S1b VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 VPWR S0 S0b VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 VPWR xb X VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux4_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs1o xb S1b xlowb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNs2o xb S1 xhib VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 VGND S1 S1b VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 VGND S0 S0b VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN4 VGND xb X VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs1o xb S1 xlowb VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPs2o xb S1b xhib VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 VPWR S1 S1b VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 VPWR S0 S0b VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 VPWR xb X VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux4_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNs1o xb S1b xlowb VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNs2o xb S1 xhib VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN1 VGND S1 S1b VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 VGND S0 S0b VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN4 VGND xb X VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPs1o xb S1 xlowb VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPs2o xb S1b xhib VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP1 VPWR S1 S1b VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP2 VPWR S0 S0b VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP4 VPWR xb X VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__mux4_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=8 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand2_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2b_1 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nand2b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2b_2 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nand2b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand2b_4 A_N B VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand2b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3_2 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3_4 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3b_1 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nand3b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3b_2 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nand3b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand3b_4 A_N B C VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 sndB C VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand3b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4_1 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand4_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand4_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4_4 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand4_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nand4b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nand4b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand4b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nand4bb_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nand4bb_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
*.PININFO A_N:I B_N:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 Y B VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 Y C VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP3 Y D VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP0 A A_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A sndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 sndA B sndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 sndB C sndC VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN3 sndC D VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN0 A A_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nand4bb_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2_8 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=8 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=8 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor2_8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2b_1 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nor2b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2b_2 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nor2b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor2b_4 A B_N VGND VNB VPB VPWR Y
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor2b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3_1 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3_2 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3_4 A B C VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3b_1 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nor3b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3b_2 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nor3b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor3b_4 A B C_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 sndPB C Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor3b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4_1 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor4_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor4_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4_4 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor4_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nor4b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nor4b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor4b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__nor4bb_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__nor4bb_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=4 w=1.12 l=0.15
MMP3 sndPC D Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMN0 Y A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN1 Y B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN2 Y C VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMN3 Y D VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__nor4bb_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPD0 VPWR D1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 y D1 pndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPD0 VPWR D1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 y D1 pndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPD0 VPWR D1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMND0 y D1 pndC VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPD0 VPWR D1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMND0 Y D1 pndC VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPD0 VPWR D1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMND0 Y D1 pndC VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I D1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPD0 VPWR D1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNC0 pndC C1 pndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMND0 Y D1 pndC VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o2111ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o211ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ba_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ba_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21ba_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
.ENDS sky130_fd_sc_hs__o21bai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__o21bai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1_N:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMIPB1N B1 B1_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMINB1N B1 B1_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o21bai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 pndB B2 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o221ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o22ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi20 y inand nmid VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi11 sndPB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi20 y inand VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 y inand nmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi11 sndPB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi20 y inand VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi20 y inand nmid VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPaoi11 sndPB1 B2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPaoi20 y inand VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1_N:I A2_N:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi10 nmid B1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi11 nmid B2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMPnand0 inand A1_N VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPnand1 inand A2_N VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__o2bb2ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPC0 VPWR C1 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNC0 y C1 pndB VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I C1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPC0 VPWR C1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 pndB B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNC0 Y C1 pndB VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o311ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o31ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPA2 sndA2 A3 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPB1 sndB1 B2 y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB1 y B2 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 sndA2 A3 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 sndB1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB1 sndB1 B2 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB1 Y B2 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o32ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA3 sndA3 A4 y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41a_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA3 sndA3 A4 y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41a_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA3 sndA3 A4 y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 y VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIPX X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNB0 y B1 pndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMINX X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41a_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPA3 sndA3 A4 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41ai_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPA3 sndA3 A4 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41ai_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
*.PININFO A1:I A2:I A3:I A4:I B1:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMPA0 VPWR A1 sndA1 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPA3 sndA3 A4 Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPB0 VPWR B1 Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMNA0 pndA A1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA1 pndA A2 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA2 pndA A3 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNA3 pndA A4 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNB0 Y B1 pndA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__o41ai_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=0.84 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2b_1 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2b_2 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or2b_4 A B_N VGND VNB VPB VPWR X
*.PININFO A:I B_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP1 B B_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN1 B B_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or2b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3b_1 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3b_2 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or3b_4 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 sndPB C y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN3 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or3b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4_1 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4_2 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4_4 A B C D VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4b_1 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4b_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4b_2 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4b_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4b_4 A B C D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4b_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4bb_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=1 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4bb_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I D_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP1 sndPA B sndPB VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP2 sndPB C sndPC VPB pfet_01v8 m=2 w=1.0 l=0.15
MMP3 sndPC D y VPB pfet_01v8 m=2 w=1.0 l=0.15
MMIP2 C C_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP3 D D_N VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMIP4 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN1 y B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN2 y C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMN3 y D VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMIN2 C C_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN3 D D_N VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIN4 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__or4bb_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
MI98 net105 D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 net105 SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net176 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net213 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI677 M1 RESET net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net160 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net160 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net145 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net145 net117 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net117 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 net213 net117 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI42 net105 clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net125 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net125 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net117 RESET net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net117 S0 net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net116 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 net105 D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 net105 sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net265 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net213 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI9 net117 S0 net268 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net265 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net216 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net257 net117 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net257 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net117 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net268 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net241 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 net105 clkpos M0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI656 M0 clkneg net241 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net216 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net213 net117 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI661 Q_N net117 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfbbn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
MI98 net105 D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 net105 SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net176 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net213 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI677 M1 RESET net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net160 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net160 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net145 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net145 net117 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net117 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI652 net213 net117 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI42 net105 clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net125 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net125 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net117 RESET net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net117 S0 net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net116 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 net105 D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 net105 sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net265 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net213 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI9 net117 S0 net268 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net265 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net216 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net257 net117 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net257 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net117 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net268 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net241 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 net105 clkpos M0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI656 M0 clkneg net241 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net216 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net213 net117 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI661 Q_N net117 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfbbn_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I
*.PININFO VPWR:I Q:O Q_N:O
MI98 net105 D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 net105 SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 RESET RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI676 M1 M0 net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI675 net176 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net213 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI677 M1 RESET net176 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI648 M0 clkpos net153 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 net153 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 S0 clkneg net145 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net145 net117 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N net117 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 net213 net117 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI42 net105 clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI668 S0 clkpos net128 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI667 net128 M1 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI630 net117 RESET net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI3 net117 S0 net116 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI7 net116 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 net105 D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 net105 sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI679 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI669 S0 clkneg net265 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net213 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI9 net117 S0 net268 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI670 net265 M1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI678 net216 RESET VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI662 net257 net117 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 S0 clkpos net257 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI10 net117 SET_B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI11 net268 RESET VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 net241 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 net105 clkpos M0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI656 M0 clkneg net241 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI643 RESET RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI680 M1 M0 net216 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI663 net213 net117 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI661 Q_N net117 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfbbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O Q_N:O
MI642 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI651 Q_N s0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net94 s0 net128 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net128 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net109 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net109 M1 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net104 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net189 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net189 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net104 net94 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI666 net148 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net148 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net148 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net217 net94 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net94 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net217 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net94 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net196 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net196 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net189 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net189 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI661 Q_N s0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O Q_N:O
MI642 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI651 Q_N s0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net92 s0 net126 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net126 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net119 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net107 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net107 M1 net119 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net91 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net187 s0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI653 Q net187 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI654 net91 net92 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI666 net146 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net146 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net146 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net215 net92 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net92 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net215 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net92 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net194 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net194 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net187 s0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net187 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI661 Q_N s0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI642 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net87 s0 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net114 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net102 M1 net114 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net97 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net174 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net174 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net97 net87 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI666 net137 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net202 net87 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net87 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net202 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net87 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net181 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net181 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net174 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net174 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrtn_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI642 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net87 s0 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net114 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net102 M1 net114 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net86 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net174 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI653 Q net174 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI654 net86 net87 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI666 net137 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net202 net87 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net87 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net202 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net87 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net181 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net181 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net174 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net174 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI642 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net87 s0 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net114 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net102 M1 net114 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net86 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net174 s0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI653 Q net174 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI654 net86 net87 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI666 net137 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net202 net87 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net87 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net202 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net87 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net181 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net181 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net174 s0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net174 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI642 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net87 s0 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI33 net114 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI4 M0 clkpos net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net102 M1 net114 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 s0 clkneg net97 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net174 s0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 Q net174 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI654 net97 net87 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI666 net137 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI635 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net202 net87 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net87 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 s0 clkpos net202 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 net87 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI30 net181 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI31 M0 clkneg net181 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI663 net174 s0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI660 Q net174 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfrtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI662 net159 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net159 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net138 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI669 S0 clkpos net138 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI661 Q_N S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI663 net199 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI660 Q net199 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net98 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net98 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI27 net243 S1 net215 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI34 S0 clkpos net187 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI657 net227 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI653 Q net199 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI644 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI25 net215 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI651 Q_N S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkpos net206 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI652 net199 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI656 M1 M0 net227 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net206 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI36 net187 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI26 S0 clkneg net243 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sdfsbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI645 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI663 net195 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net195 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net130 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net130 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net122 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI669 S0 clkpos net122 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net107 VPB pfet_01v8 m=2 w=0.84 l=0.15
MI37 net107 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI661 Q_N S0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 S0 clkpos net219 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI27 net239 S1 net187 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net230 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net199 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net230 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI36 net219 M0 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI26 S0 clkneg net239 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net199 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net195 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI644 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI25 net187 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI653 Q net195 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI651 Q_N S0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__sdfsbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI645 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI663 net165 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 Q net165 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net104 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net104 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net96 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI669 S0 clkpos net96 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net84 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI37 net84 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI34 S0 clkpos net189 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI27 net209 S1 net157 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net200 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net169 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net200 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI36 net189 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI26 S0 clkneg net209 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net169 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net165 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI644 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI25 net157 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI653 Q net165 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sdfstp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI645 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI663 net165 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI660 Q net165 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net109 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net109 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net96 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI669 S0 clkpos net96 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net84 VPB pfet_01v8 m=2 w=0.84 l=0.15
MI37 net84 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI34 S0 clkpos net212 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI27 net209 S1 net157 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net200 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net169 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net200 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI36 net212 M0 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI26 S0 clkneg net209 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net169 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net165 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI644 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI25 net157 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI653 Q net165 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sdfstp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I SET_B:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI645 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI47 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI663 net165 S0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI660 Q net165 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI659 M1 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI662 net104 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkneg net104 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI6 net96 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI669 S0 clkpos net96 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI24 S0 SET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI648 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI38 S0 clkneg net84 VPB pfet_01v8 m=2 w=0.84 l=0.15
MI37 net84 M0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI45 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI34 S0 clkpos net189 VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI27 net209 S1 net157 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI647 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI655 M0 clkpos net200 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 M1 M0 net196 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net200 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI36 net189 M0 VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MI26 S0 clkneg net209 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI46 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI657 net196 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 net165 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI644 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI25 net157 SET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI653 Q net165 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sdfstp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net129 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net129 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net120 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net120 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI661 Q_N net153 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI662 net153 S1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI644 S0 clkpos net177 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 net189 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI660 Q_N net153 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net177 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI659 M0 clkneg net189 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI647 net153 S1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__sdfxbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O Q_N:O
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net132 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net132 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net120 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net120 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI661 Q_N net153 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI662 net153 S1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI644 S0 clkpos net196 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 net160 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI660 Q_N net153 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI643 net196 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI659 M0 clkneg net160 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI647 net153 S1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
.ENDS sky130_fd_sc_hs__sdfxbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net75 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net75 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net54 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 S0 clkneg net54 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 net122 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 net138 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI659 M0 clkneg net138 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net122 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfxtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net78 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net78 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net71 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 S0 clkneg net71 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 net163 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 net155 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI659 M0 clkneg net155 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI644 S0 clkpos net163 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfxtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI652 M1 clkpos S0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI649 S1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI639 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net78 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI656 net78 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI641 net54 S1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S1 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI642 S0 clkneg net54 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI103 n1 SCD VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI104 n0 sceb VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI643 net163 S1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI640 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI658 net155 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S1 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI653 M1 clkneg S0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI659 M0 clkneg net155 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 S1 S0 VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MI644 S0 clkpos net163 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__sdfxtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net88 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net88 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net76 CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI658 net76 m1 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI22 net63 SCE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI21 net116 GATE net63 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net76 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI43 net116 clkneg M0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI42 net116 clkpos M0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net123 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net123 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI24 net116 SCE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI657 net112 CLK VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI656 net76 m1 net112 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI23 net116 GATE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net76 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__sdlclkp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net88 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net88 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net76 CLK VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI658 net76 m1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI22 net63 SCE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI21 net116 GATE net63 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net76 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI43 net116 clkneg M0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI42 net116 clkpos M0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net123 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net123 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI24 net116 SCE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI657 net112 CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net76 m1 net112 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI23 net116 GATE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net76 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__sdlclkp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
*.PININFO CLK:I GATE:I SCE:I VGND:I VNB:I VPB:I VPWR:I GCLK:O
MI662 net88 m1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI664 M0 clkpos net88 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 net76 CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net76 m1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 m1 M0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI22 net63 SCE VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI21 net116 GATE net63 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI45 clkpos CLK VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI660 GCLK net76 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI43 net116 clkneg M0 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI42 net116 clkpos M0 VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI20 m1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI655 M0 clkneg net123 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI654 net123 m1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI24 net116 SCE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI657 net112 CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net76 m1 net112 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI23 net116 GATE VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MI46 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI44 clkpos CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI653 GCLK net76 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__sdlclkp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI14 net154 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net154 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net143 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net126 q1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net126 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI660 Q_N q1 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI659 M0 clkneg net143 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 q1 S0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI33 net111 deneg VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 net102 sceneg db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI46 VPWR SCD net102 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI31 net99 D net111 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI42 net99 SCE db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI40 net82 q1 net99 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI36 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI38 VPWR DE net82 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI44 sceneg SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI661 Q_N q1 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net235 q1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net235 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net219 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net219 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI43 net99 sceneg db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 q1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI45 sceneg SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI32 net99 D net198 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net195 M1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI15 S0 clkpos net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI41 net187 q1 net99 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI39 VGND deneg net187 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI37 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net198 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI49 net166 SCE db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI48 VGND SCD net166 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sedfxbp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI14 net154 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net154 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI658 net143 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net126 q1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net126 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI660 Q_N q1 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI659 M0 clkneg net143 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 q1 S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI33 net111 deneg VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 net107 sceneg db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI46 VPWR SCD net107 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI31 net99 D net111 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI42 net99 SCE db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI40 net91 q1 net99 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI36 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI38 VPWR DE net91 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI44 sceneg SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI661 Q_N q1 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI641 net235 q1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net235 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI656 net214 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net214 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI43 net99 sceneg db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 q1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI45 sceneg SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI32 net99 D net175 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net195 M1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI15 S0 clkpos net195 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI41 net182 q1 net99 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI39 VGND deneg net182 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI37 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net175 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI49 net166 SCE db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI48 VGND SCD net166 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sedfxbp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI14 net146 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net146 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI658 net135 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net118 q1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net118 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 M0 clkneg net135 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 q1 S0 VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI33 net107 deneg VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 net98 sceneg db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI46 VPWR SCD net98 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI31 net95 D net107 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI42 net95 SCE db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI40 net78 q1 net95 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI36 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI38 VPWR DE net78 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI44 sceneg SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net227 q1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net227 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI656 net211 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net211 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI43 net95 sceneg db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 q1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI45 sceneg SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI32 net95 D net190 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net187 M1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI15 S0 clkpos net187 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI41 net179 q1 net95 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI39 VGND deneg net179 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI37 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net190 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI49 net158 SCE db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI48 VGND SCD net158 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sedfxtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI14 net146 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net146 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI658 net114 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net118 q1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net118 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 M0 clkneg net114 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 q1 S0 VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI33 net107 deneg VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 net98 sceneg db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI46 VPWR SCD net98 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI31 net95 D net107 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI42 net95 SCE db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI40 net78 q1 net95 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI36 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI38 VPWR DE net78 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI44 sceneg SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net222 q1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net222 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI656 net211 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net211 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI43 net95 sceneg db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 q1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI45 sceneg SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI32 net95 D net190 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net187 M1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI15 S0 clkpos net187 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI41 net179 q1 net95 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI39 VGND deneg net179 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI37 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net190 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI49 net163 SCE db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI48 VGND SCD net163 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sedfxtp_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI14 net146 M1 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI637 clkpos clkneg VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI13 S0 clkneg net146 VPB pfet_01v8 m=1 w=1.0 l=0.15
MI651 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI645 Q S0 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI658 net135 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI638 clkneg CLK VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI643 net118 q1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.15
MI639 M1 M0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MI644 S0 clkpos net118 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI659 M0 clkneg net135 VPB pfet_01v8 m=1 w=0.42 l=0.15
MI17 q1 S0 VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI33 net107 deneg VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI47 net98 sceneg db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI46 VPWR SCD net98 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI31 net95 D net107 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI42 net95 SCE db VPB pfet_01v8 m=1 w=0.64 l=0.15
MI40 net78 q1 net95 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI36 deneg DE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI38 VPWR DE net78 VPB pfet_01v8 m=1 w=0.64 l=0.15
MI44 sceneg SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI634 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI636 clkpos clkneg VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI635 clkneg CLK VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI641 net227 q1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI642 S0 clkneg net227 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI648 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI646 Q S0 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI656 net211 M1 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI657 M0 clkpos net211 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI43 net95 sceneg db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI18 q1 S0 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI45 sceneg SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI32 net95 D net190 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI16 net187 M1 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI15 S0 clkpos net187 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI41 net179 q1 net95 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI39 VGND deneg net179 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI37 deneg DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI34 net190 DE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI49 net158 SCE db VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI48 VGND SCD net158 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
.ENDS sky130_fd_sc_hs__sedfxtp_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor2_1 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnand1 sndNA B inand VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 nmid A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 nmid B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPnand0 inand A VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPnand1 inand B VPWR VPB pfet_01v8 m=1 w=0.84 l=0.15
MMPaoi10 VPWR A sndPA VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi11 sndPA B Y VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xnor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor2_2 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNnand1 sndNA B inand VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi10 nmid A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi11 nmid B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPnand0 inand A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnand1 inand B VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 VPWR A sndPA VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi11 sndPA B Y VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xnor2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor2_4 A B VGND VNB VPB VPWR Y
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNnand0 VGND A sndNA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNnand1 sndNA B inand VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMNaoi10 nmid A VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi11 nmid B VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi20 Y inand nmid VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMPnand0 inand A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPnand1 inand B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMPaoi10 VPWR A sndPA VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi11 sndPA B Y VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi20 Y inand VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xnor2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN3 X net57 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 mid1 Cb net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI2 mid2 C net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP3 X net57 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 mid1 C net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI7 mid2 Cb net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__xnor3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN3 X net57 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 mid1 Cb net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI2 mid2 C net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP3 X net57 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI650 mid1 C net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI7 mid2 Cb net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__xnor3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xnor3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN3 X net57 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI649 mid1 Cb net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI2 mid2 C net57 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMIP3 X net57 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI650 mid1 C net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI7 mid2 Cb net57 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
.ENDS sky130_fd_sc_hs__xnor3_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNnor0 inor A VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNnor1 inor B VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15
MMNaoi10 VGND A sndNA VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi11 sndNA B X VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMNaoi20 X inor VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPnor0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA B inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid A VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi11 pmid B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MMPaoi20 X inor pmid VPB pfet_01v8 m=1 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor2_2 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNnor0 inor A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNnor1 inor B VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MMNaoi10 VGND A sndNA VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi11 sndNA B X VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi20 X inor VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MMPnor0 VPWR A sndPA VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPnor1 sndPA B inor VPB pfet_01v8 m=1 w=1.0 l=0.15
MMPaoi10 pmid A VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi11 pmid B VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMPaoi20 X inor pmid VPB pfet_01v8 m=2 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xor2_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor2_4 A B VGND VNB VPB VPWR X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNnor0 inor A VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNnor1 inor B VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMNaoi10 VGND A sndNA VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi11 sndNA B X VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MMNaoi20 X inor VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MMPnor0 VPWR A sndPA VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPnor1 sndPA B inor VPB pfet_01v8 m=2 w=1.0 l=0.15
MMPaoi10 pmid A VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi11 pmid B VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMPaoi20 X inor pmid VPB pfet_01v8 m=4 w=1.12 l=0.15
.ENDS sky130_fd_sc_hs__xor2_4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor3_1 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIP3 X net117 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI650 mid1 Cb net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 mid2 C net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIN3 X net117 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 mid1 C net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 mid2 Cb net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__xor3_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIP3 X net117 VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MI650 mid1 Cb net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 mid2 C net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIN3 X net117 VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 mid1 C net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 mid2 Cb net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__xor3_2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hs__xor3_4 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIP3 X net117 VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MI650 mid1 Cb net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI1 mid2 C net117 VPB pfet_01v8 m=1 w=0.84 l=0.15
MI33 Cb C VPWR VPB pfet_01v8 m=1 w=0.64 l=0.15
MI45 Ab A VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI47 Abb Ab VPWR VPB pfet_01v8 m=1 w=1.0 l=0.15
MI19 mid1 Bb Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MI16 Bb B VPWR VPB pfet_01v8 m=1 w=1.12 l=0.15
MI23 mid1 B Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI26 mid2 Bb Abb VPB pfet_01v8 m=1 w=0.64 l=0.15
MI27 mid2 B Ab VPB pfet_01v8 m=1 w=0.84 l=0.15
MMIN3 X net117 VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
MI34 Cb C VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI649 mid1 C net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI2 mid2 Cb net117 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI44 Ab A VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI46 Abb Ab VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI17 Bb B VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15
MI24 Ab B mid1 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI25 Abb Bb mid1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15
MI28 Abb B mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
MI29 Ab Bb mid2 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15
.ENDS sky130_fd_sc_hs__xor3_4
